module MPDataLoader (
    input clk,
    input rst
);
    
    always @ (*) begin
    end

    always @ (posedge clk) begin
        if (rst) begin
        end
        else begin
        end
    end
endmodule