module CVDataLoader (
    
);
    
endmodule
