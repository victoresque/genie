module CVCore (
    
);
    
endmodule
